// Copyright (C) 2016  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
// Created on Sun Oct 20 21:13:50 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module HW6P2 (
    reset,clock,A,B,C,D,PBGNT,MACK,CONT,
    PBREQ,CNTLD,CMREQ,CLD,CE);

    input reset;
    input clock;
    input A;
    input B;
    input C;
    input D;
    input PBGNT;
    input MACK;
    input CONT;
    tri0 reset;
    tri0 A;
    tri0 B;
    tri0 C;
    tri0 D;
    tri0 PBGNT;
    tri0 MACK;
    tri0 CONT;
    output PBREQ;
    output CNTLD;
    output CMREQ;
    output CLD;
    output CE;
    reg PBREQ;
    reg CNTLD;
    reg CMREQ;
    reg CLD;
    reg CE;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3,S4=4,S5=5;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or A or B or C or D or PBGNT or MACK or CONT)
    begin
        if (reset) begin
            reg_fstate <= S0;
            PBREQ <= 1'b0;
            CNTLD <= 1'b0;
            CMREQ <= 1'b0;
            CLD <= 1'b0;
            CE <= 1'b0;
        end
        else begin
            PBREQ <= 1'b0;
            CNTLD <= 1'b0;
            CMREQ <= 1'b0;
            CLD <= 1'b0;
            CE <= 1'b0;
            case (fstate)
                S0: begin
                    if ((((~(A) & ~(B)) & ~(C)) & ~(D)))
                        reg_fstate <= S0;
                    else if ((((A | B) | C) | D))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;
                end
                S1: begin
                    if (~(PBGNT))
                        reg_fstate <= S1;
                    else if (PBGNT)
                        reg_fstate <= S2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;

                    PBREQ <= 1'b1;
                end
                S2: begin
                    if (~(MACK))
                        reg_fstate <= S2;
                    else if (MACK)
                        reg_fstate <= S3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;

                    CMREQ <= 1'b1;

                    CNTLD <= 1'b1;
                end
                S3: begin
                    reg_fstate <= S4;

                    CE <= 1'b1;
                end
                S4: begin
                    if (~(CONT))
                        reg_fstate <= S0;
                    else if (CONT)
                        reg_fstate <= S5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S4;

                    CLD <= 1'b1;
                end
                S5: begin
                    if (~(MACK))
                        reg_fstate <= S5;
                    else if (MACK)
                        reg_fstate <= S3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S5;

                    CMREQ <= 1'b1;
                end
                default: begin
                    PBREQ <= 1'bx;
                    CNTLD <= 1'bx;
                    CMREQ <= 1'bx;
                    CLD <= 1'bx;
                    CE <= 1'bx;
                    $display ("%d: Reach undefined state", $time);
                end
            endcase
        end
    end
endmodule // HW6P2
