library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cc is 
port ( clk : in std_logic;
		 compin, reset: in std_logic;
		 Q3 : out std_logic );
end entity CC:

architecture behavioral of CC is
begin
	process(clk, reset)
	begin
		
		



end
